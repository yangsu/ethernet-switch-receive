--LIBRARY ieee;
--USE ieee.std_logic_1164.all;
--USE ieee.numeric_std.all;
--
--ENTITY receive IS
--	PORT (
--		aclr				:	IN 	STD_LOGIC;
--		clk25				:	IN STD_LOGIC;
--		clk50				:	IN STD_LOGIC;
--		data_in				:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--		data_in_valid		: 	IN STD_LOGIC;
--		hold				: 	IN STD_LOGIC;
--	);
--END receive;
--
--	COMPONENT inputProcessor IS
--		PORT (	aclr			:	IN STD_LOGIC;
--				clk25			:	IN STD_LOGIC;
--				clk50			:	IN STD_LOGIC;
--				data_in			:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
--				data_in_valid	: 	IN STD_LOGIC;
--				data_out		:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
--				data_out_valid	:	OUT STD_LOGIC;
--				crc				:	OUT STD_LOGIC;
--				frame_length	:	OUT STD_LOGIC_VECTOR(11 DOWNTO 0); -- Max frame size is 1542 bytes
--				receive_state	:	OUT STD_LOGIC;
--				hold_state		:	OUT STD_LOGIC;
--				reset_state		:	OUT STD_LOGIC);
--	END COMPONENT;
--
--ARCHITECTURE rcv OF receive IS
--
--END rcv